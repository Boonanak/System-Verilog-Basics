module tb;
    hello_world hw();
endmodule